module detection_unit(
    input [3:0] curr_rs, curr_rt,
    input [3:0] d_rd, e_rd,
    input branch,
    output hazard_sig,

);







endmodule