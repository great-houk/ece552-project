//////////////////////////////////////
//
// Memory -- single cycle version
//
// written for CS/ECE 552, Spring '07
// Pratap Ramamurthy, 19 Mar 2006
//
// Modified for CS/ECE 552, Spring '18
// Gokul Ravi, 08 Mar 2018
//
// This is a byte-addressable,
// 16-bit wide memory
// Note: The last bit of the address has to be 0.
//
// All reads happen combinationally with zero delay.
// All writes occur on rising clock edge.
// Concurrent read and write not allowed.
//
// On reset, memory loads from file "loadfile_all.img".
// (You may change the name of the file in
// the $readmemh statement below.)
// File format:
//     @0
//     <hex data 0>
//     <hex data 1>
//     ...etc
//
//
//////////////////////////////////////

module memory1c_instr (data_out, data_in, addr, enable, wr, clk, rst);

   parameter ADDR_WIDTH = 16;
   output  [15:0] data_out;
   input [15:0]   data_in;
   input [ADDR_WIDTH-1 :0]   addr;
   input          enable;
   input          wr;
   input          clk;
   input          rst;
   wire [15:0]    data_out;
   
   reg [15:0]      mem [0:2**ADDR_WIDTH-1];
   reg            loaded;
   
   // TODO: Fix this
   wire [15:0] mem_read_data;
   assign mem_read_data = mem[addr[ADDR_WIDTH-1 :1]];
   assign data_out = (enable & (~wr))? {mem[addr[ADDR_WIDTH-1 :1]]}: 0;
   initial begin
      loaded = 0;
   end

   always @(posedge clk) begin
      if (rst) begin
         //load program.img
         if (!loaded) begin
            $readmemh("program.img", mem);
            loaded = 1;
         end
          
      end
      else begin
         if (enable & wr) begin
	        mem[addr[ADDR_WIDTH-1 :1]] = data_in[15:0];       // The actual write
         end
      end
   end
endmodule



module memory1c (data_out, data_in, addr, enable, wr, clk, rst);

   parameter ADDR_WIDTH = 16;
   output  [15:0] data_out;
   input [15:0]   data_in;
   input [ADDR_WIDTH-1 :0]   addr;
   input          enable;
   input          wr;
   input          clk;
   input          rst;
   wire [15:0]    data_out;
   
   reg [15:0]      mem [0:2**ADDR_WIDTH-1];
   reg            loaded;
   
   // TODO: Fix this
   wire [15:0] mem_read_data;
   assign mem_read_data = mem[addr[ADDR_WIDTH-1 :1]];
   assign data_out = (enable & (~wr))? {mem[addr[ADDR_WIDTH-1 :1]]}: 0;
   initial begin
      loaded = 0;
   end

	integer i;
   always @(posedge clk) begin
      if (rst) begin
         //load loadfile_all.img
        //  if (!loaded) begin
        //     $readmemh("loadfile_all_data.img", mem);
        //     loaded = 1;
        //  end
		
		// Set the memory to 0 on reset
		for (i = 0; i < 2**ADDR_WIDTH; i = i + 1) begin
			mem[i] = 16'h0000;
		end
		loaded = 1;  
      end
      else begin
         if (enable & wr) begin
	        mem[addr[ADDR_WIDTH-1 :1]] = data_in[15:0];       // The actual write
         end
      end
   end


endmodule 
