module forwarding_unit(
	input clk, rst_n,
	input ex_ex_forwarding,
	input ex_mem_forwarding,
	input mem_mem_forwarding,
	input [15:0] m_alu_result,
	input 
);

endmodule